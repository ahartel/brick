
package clk_period;
	int period = 6;
endpackage
